--- !ruby/object:Hangman
file: 5desk.txt
tries: 6
max_tries: 10
guessed:
- l
- m
- e
- s
word: slimmer
